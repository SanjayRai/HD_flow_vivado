/*
------------------------------------------------------------------
--      _____
--     /     \
--    /____   \____
--   / \===\   \==/
--  /___\===\___\/  AVNET
--       \======/
--        \====/    
------------------------------------------------------------------
--
-- This design is the property of Avnet.  Publication of this
-- design is not authorized without written consent from Avnet.
-- 
-- Please direct any questions to:  technical.support@avnet.com
--
-- Disclaimer:
--    Avnet, Inc. makes no warranty for the use of this code or design.
--    This code is provided  "As Is". Avnet, Inc assumes no responsibility for
--    any errors, which may appear in this code, nor does it make a commitment
--    to update the information contained herein. Avnet, Inc specifically
--    disclaims any implied warranties of fitness for a particular purpose.
--                     Copyright(c) 2010 Avnet, Inc.
--                             All rights reserved.
--
------------------------------------------------------------------
--
-- Create Date:         Jan 20, 2010
-- Design Name:         DVI_Pass_Through_Demo
-- Module Name:         PB_FMC_DVIDP_CONFIG
-- Project Name:        DVI_Pass_Through_Demo
-- Target Devices:      Spartan-6
-- Avnet Boards:        FMC-DVI/DP
--
-- Tool versions:       ISE 12.2
--
-- Description:         This is a module for storing a program for the KCPSM3 (aka Pico-Blaze)
--                      The code is assembled as "pbt3" (should be pbt3 for spartan 3)
--
--                      Ingredients: 1 18kb Block Ram
--
-- Dependencies:        
--
-- Revision:            Jan 20, 2010: 1.00 Initial Version
--                      Sep 07, 2010: 1.01 Update for 12.2
--
------------------------------------------------------------------
*/

module PB_FMC_DVIDP_CONFIG(
	CLK, ADDRESS, INSTRUCTION,
	LOAD_CLK, LOAD_ADDRESS, LOAD_INSTRUCTION, LOAD_WE
	);

input			CLK;
input	[9:0]	ADDRESS;
output	[17:0]	INSTRUCTION;

// Load interface for reloading program
input			LOAD_CLK;
input	[9:0]	LOAD_ADDRESS;
input	[17:0]	LOAD_INSTRUCTION;
input			LOAD_WE;

RAMB16_S18_S18	#(
      .INIT_00(256'h4003400F002F002600200013400F400A1400A01C40025002A008400300134005),
      .INIT_01(256'hA00000C80A64C000000000C80A64C000000100C80A64C00000004002540FA008),	
      .INIT_02(256'h0070A000003806040502003806F10506E0110040A000003806040504E01100E0),	
      .INIT_03(256'h007485011850B40029010074681100A0A00000380610050A003806B30508E011),	
      .INIT_04(256'h1870B4002901007485011850B40029010074681100A0A00000791860B4002901),	
      .INIT_05(256'h601000746812B00040006010B40029010074681100A0A00000791860B4000074),	
      .INIT_06(256'h407C08FF0900A0000074C801681100A0B40029010055A00000746813B0004001),	
      .INIT_07(256'h000000010806010840B1007C090140B1B0002901007C090140B1007C08FF0901),	
      .INIT_08(256'h547DC10100BE0A05C0010008D800A001400100BE0A0AC001000C00BE0A05C001),	
      .INIT_09(256'hA00000BE0A05C0010008490100BE0A0AC001000C00BE0A05C001C002A0011090),	
      .INIT_0A(256'h00BE0A05C001000800BE0A05C001000200BE0A05C001000C00BE0A05C0010003),	
      .INIT_0B(256'hCB060B0CA00000BE0A05C001000300BE0A05C001000C00BE0A05C0010002A000),	
      .INIT_0C(256'h00BE0AFA00BE0AFA00BE0AFA00BE0AFAA00054BECA0154C3CB02CB0150C32B01),	
      .INIT_0D(256'h0000000000000000000000000000000000000000000000008000A00054C8C001),	
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_3F(256'h40D3000000000000000000000000000000000000000000000000000000000000),
      .INITP_00(256'h88F39CF0C2C39EC93249CECB2749CEC9D273B0C22C308B08B232323C3FFF030F),
      .INITP_01(256'h0000000000000000000000EDCCCCB75D4B232322C8C8C8C8B20C8C80DC803232),
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INITP_07(256'hC000000000000000000000000000000000000000000000000000000000000000))
rom(	
	// Port A: Read Port
	.CLKA(CLK), .ADDRA(ADDRESS),
	.DIA(16'h0000), .DIPA(2'b00), .WEA(1'b0),
	.DOA(INSTRUCTION[15:0]), .DOPA(INSTRUCTION[17:16]),
	.ENA(1'b1), .SSRA(1'b0),
	// port B: Load (write) port
	.CLKB(LOAD_CLK), .ADDRB(LOAD_ADDRESS), 
	.DIB(LOAD_INSTRUCTION[15:0]), .DIPB(LOAD_INSTRUCTION[17:16]), .WEB(LOAD_WE),
	.DOB(), .DOPB(),
	.ENB(1'b1), .SSRB(1'b0)
	);


endmodule
